magic
tech sky130A
magscale 1 2
timestamp 1701930086
<< metal3 >>
rect -406 812 406 840
rect -406 -812 322 812
rect 386 -812 406 812
rect -406 -840 406 -812
<< via3 >>
rect 322 -812 386 812
<< mimcap >>
rect -366 760 74 800
rect -366 -760 -326 760
rect 34 -760 74 760
rect -366 -800 74 -760
<< mimcapcontact >>
rect -326 -760 34 760
<< metal4 >>
rect 306 812 402 828
rect -327 760 35 761
rect -327 -760 -326 760
rect 34 -760 35 760
rect -327 -761 35 -760
rect 306 -812 322 812
rect 386 -812 402 812
rect 306 -828 402 -812
<< properties >>
string FIXED_BBOX -406 -840 114 840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.20 l 8.00 val 39.076 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
