magic
tech sky130A
magscale 1 2
timestamp 1701909091
<< error_p >>
rect -29 281 29 287
rect -29 247 -17 281
rect -29 241 29 247
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect -29 -287 29 -281
<< nwell >>
rect -220 -419 220 419
<< pmos >>
rect -24 -200 24 200
<< pdiff >>
rect -82 188 -24 200
rect -82 -188 -70 188
rect -36 -188 -24 188
rect -82 -200 -24 -188
rect 24 188 82 200
rect 24 -188 36 188
rect 70 -188 82 188
rect 24 -200 82 -188
<< pdiffc >>
rect -70 -188 -36 188
rect 36 -188 70 188
<< nsubdiff >>
rect -184 349 -88 383
rect 88 349 184 383
rect -184 287 -150 349
rect 150 287 184 349
rect -184 -349 -150 -287
rect 150 -349 184 -287
rect -184 -383 -88 -349
rect 88 -383 184 -349
<< nsubdiffcont >>
rect -88 349 88 383
rect -184 -287 -150 287
rect 150 -287 184 287
rect -88 -383 88 -349
<< poly >>
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect -24 200 24 231
rect -24 -231 24 -200
rect -33 -247 33 -231
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -297 33 -281
<< polycont >>
rect -17 247 17 281
rect -17 -281 17 -247
<< locali >>
rect -184 349 -88 383
rect 88 349 184 383
rect -184 287 -150 349
rect 150 287 184 349
rect -33 247 -17 281
rect 17 247 33 281
rect -70 188 -36 204
rect -70 -204 -36 -188
rect 36 188 70 204
rect 36 -204 70 -188
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -184 -349 -150 -287
rect 150 -349 184 -287
rect -184 -383 -88 -349
rect 88 -383 184 -349
<< viali >>
rect -17 247 17 281
rect -70 -188 -36 188
rect 36 -188 70 188
rect -17 -281 17 -247
<< metal1 >>
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect -76 188 -30 200
rect -76 -188 -70 188
rect -36 -188 -30 188
rect -76 -200 -30 -188
rect 30 188 76 200
rect 30 -188 36 188
rect 70 -188 76 188
rect 30 -200 76 -188
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect 17 -281 29 -247
rect -29 -287 29 -281
<< properties >>
string FIXED_BBOX -167 -366 167 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.24 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
