magic
tech sky130A
timestamp 1701909091
<< nmos >>
rect -12 -50 12 50
<< ndiff >>
rect -41 44 -12 50
rect -41 -44 -35 44
rect -18 -44 -12 44
rect -41 -50 -12 -44
rect 12 44 41 50
rect 12 -44 18 44
rect 35 -44 41 44
rect 12 -50 41 -44
<< ndiffc >>
rect -35 -44 -18 44
rect 18 -44 35 44
<< poly >>
rect -12 50 12 63
rect -12 -63 12 -50
<< locali >>
rect -35 44 -18 52
rect -35 -52 -18 -44
rect 18 44 35 52
rect 18 -52 35 -44
<< viali >>
rect -35 -44 -18 44
rect 18 -44 35 44
<< metal1 >>
rect -38 44 -15 50
rect -38 -44 -35 44
rect -18 -44 -15 44
rect -38 -50 -15 -44
rect 15 44 38 50
rect 15 -44 18 44
rect 35 -44 38 44
rect 15 -50 38 -44
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.24 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
