magic
tech sky130A
magscale 1 2
timestamp 1701930086
<< metal3 >>
rect -396 412 396 440
rect -396 -412 312 412
rect 376 -412 396 412
rect -396 -440 396 -412
<< via3 >>
rect 312 -412 376 412
<< mimcap >>
rect -356 360 64 400
rect -356 -360 -316 360
rect 24 -360 64 360
rect -356 -400 64 -360
<< mimcapcontact >>
rect -316 -360 24 360
<< metal4 >>
rect 296 412 392 428
rect -317 360 25 361
rect -317 -360 -316 360
rect 24 -360 25 360
rect -317 -361 25 -360
rect 296 -412 312 412
rect 376 -412 392 412
rect 296 -428 392 -412
<< properties >>
string FIXED_BBOX -396 -440 104 440
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.10 l 4.00 val 19.118 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
